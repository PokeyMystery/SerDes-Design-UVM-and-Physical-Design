`include"interface.sv"
`include "seq_item.sv"
//`include "base_seq.sv"
`include "sequencer.sv"
`include "driver.sv"

`include "monitor.sv"
//`include "subscriber.sv"

`include "scb.sv"
`include "agent.sv"
`include "env.sv"


